-- ---------------------------------------------------------------------
-- @file : bench.vhd testbench for the EP4CE6 OMDAZZ Board
-- ---------------------------------------------------------------------
--
-- Last change: KS 14.05.2023 13:02:38
-- @project: microCore
-- @language: VHDL-93
-- @copyright (c): Klaus Schleisiek, All Rights Reserved.
-- @contributors:
--
-- @license: Do not use this file except in compliance with the License.
-- You may obtain a copy of the Public License at
-- https://github.com/microCore-VHDL/microCore/tree/master/documents
-- Software distributed under the License is distributed on an "AS IS"
-- basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.
-- See the License for the specific language governing rights and
-- limitations under the License.
--
-- @brief: General simulation test bench for microCore with RS232 umbilical
-- interface. Following ARCHITECTURE, one out of a set of constants can be
-- set to '1' in order to test specific aspects of debugger.vhd.
-- When all of the constants are set to '0', bootload_sim.vhd will be
-- executed that has been cross-compiled from bootload_sim.fs.
-- The program memory will be initialized at the start of simulation when
-- MEM_FILE := "../software/program.mem". Program.mem will be generated by
-- the cross compiler.
--
-- Version Author   Date       Changes
--  1000     ks   14-May-2023  initial version
-- ---------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE work.functions_pkg.ALL;
USE work.architecture_pkg.ALL;

ENTITY bench IS
END bench;

ARCHITECTURE testbench OF bench IS

CONSTANT prog_len   : NATURAL := 10;    -- length of sim_boot.fs
CONSTANT progload   : STD_LOGIC := '0'; -- use sim_progload.fs   progload.do   MEM_file := ""                         37 usec
CONSTANT debug      : STD_LOGIC := '0'; -- use sim_debug.fs      debug.do      MEM_FILE := "../software/program.mem"  38 usec
CONSTANT handshake  : STD_LOGIC := '0'; -- use sim_handshake.fs  handshake.do  MEM_FILE := "../software/program.mem"  60 usec
CONSTANT upload     : STD_LOGIC := '0'; -- use sim_upload.fs     upload.do     MEM_FILE := "../software/program.mem"  35 usec
CONSTANT download   : STD_LOGIC := '0'; -- use sim_download.fs   download.do   MEM_FILE := "../software/program.mem"  45 usec
CONSTANT break      : STD_LOGIC := '0'; -- use sim_break.fs      break.do      MEM_FILE := "../software/program.mem" 210 usec

COMPONENT fpga PORT (                        -- pins
   reset_n     : IN    STD_LOGIC;             --  25
   clock       : IN    STD_LOGIC;             --  23  external clock input
-- Demoboard specific pins                    
   keys_n      : IN    UNSIGNED(3 DOWNTO 0);  --  91, 90, 89, 88 <= used as interrupt input during simulation
   beep        : OUT   STD_LOGIC;             -- 110
   leds_n      : OUT   UNSIGNED(3 DOWNTO 0);  --  84, 85, 86, 87
-- temp sensor                                
   SCL         : OUT   STD_LOGIC;             -- 112
   SDA         : INOUT STD_LOGIC;             -- 113
-- serial E2prom                              
   I2C_SCL     : OUT   STD_LOGIC;             --  99
   I2C_SDA     : INOUT STD_LOGIC;             --  98
-- IR es ist mir unklar, ob das ein Sender oder ein Empf�nger ist, deshal erstmal auskommentiert
--   IR          : ????? STD_LOGIC;             -- 100
-- VGA
   VGA_HSYNC   : OUT   STD_LOGIC;             -- 101
   VGA_VSYNC   : OUT   STD_LOGIC;             -- 103
   VGA_BGR     : OUT   UNSIGNED(2 DOWNTO 0);  -- 104, 105, 106
-- LCD                                        
   LCD_RS      : OUT   STD_LOGIC;             -- 141
   LCD_RW      : OUT   STD_LOGIC;             -- 138
   LCD_E       : OUT   STD_LOGIC;             -- 143
   LCD_Data    : OUT   UNSIGNED(7 DOWNTO 0);  --  11, 7, 10, 2, 3, 144, 1, 142
-- 7-Segment                                  
   DIG         : OUT   UNSIGNED(3 DOWNTO 0);  -- 137, 136, 135, 133
   SEG         : OUT   UNSIGNED(7 DOWNTO 0);  -- 127, 124, 126, 132, 129, 125, 121, 128
-- SDRAM                                      
   SD_DQ       : INOUT UNSIGNED(15 DOWNTO 0); -- 44, 46, 49, 50, 51, 52, 53, 54, 39, 38, 34, 33, 32, 31, 30, 28
   SD_A        : OUT   UNSIGNED(11 DOWNTO 0); -- 59, 75, 60, 64, 65, 66, 67, 68, 83, 80, 77, 76
   SD_BA       : OUT   UNSIGNED( 1 DOWNTO 0); -- 74, 73
   SD_LDQM     : OUT   STD_LOGIC;             -- 42
   SD_UDQM     : OUT   STD_LOGIC;             -- 55
   SD_CKE      : OUT   STD_LOGIC;             -- 58
   SD_CLK      : OUT   STD_LOGIC;             -- 43
   SD_CS_n     : OUT   STD_LOGIC;             -- 72
   SD_RAS_n    : OUT   STD_LOGIC;             -- 71
   SD_CAS_n    : OUT   STD_LOGIC;             -- 70
   SD_WE_n     : OUT   STD_LOGIC;             -- 69
-- umbilical uart for debugging
   dsu_rxd     : IN    STD_LOGIC;             -- 115  UART receive
   dsu_txd     : OUT   STD_LOGIC              -- 114  UART transmit
); END COMPONENT fpga;

SIGNAL reset_n    : STD_LOGIC;
SIGNAL xtal       : STD_LOGIC;
SIGNAL int_n      : STD_LOGIC;
SIGNAL bitout     : STD_LOGIC;

COMPONENT program_rom PORT (
   addr  : IN    program_addr;
   data  : OUT   inst_bus
); END COMPONENT;

SIGNAL debug_data   : inst_bus;
SIGNAL debug_addr   : program_addr;

SIGNAL host_rxd     : STD_LOGIC;
SIGNAL host_txd     : STD_LOGIC;
SIGNAL tx_buf       : byte;
SIGNAL send_byte    : STD_LOGIC;
SIGNAL sending      : STD_LOGIC;
SIGNAL downloading  : STD_LOGIC;
SIGNAL uploading    : STD_LOGIC;
SIGNAL host_reg     : UNSIGNED((octetts*8)-1 DOWNTO 0);
SIGNAL out_buf      : UNSIGNED((octetts*8)-1 DOWNTO 0);
SIGNAL host_buf     : byte;
SIGNAL host_full    : STD_LOGIC; -- umbilical received a data word
SIGNAL host_ack     : STD_LOGIC; -- umbilical received an ack

CONSTANT xtal_cycle : TIME := (1000000000 / xtal_frequency) * 1 ns;
CONSTANT cycle      : TIME := (1000000000 / clk_frequency) * 1 ns;
CONSTANT baud       : TIME := (cycle*clk_frequency)/umbilical_rate;
-- CONSTANT int_time   : TIME := 114260 ns + 8 * 40 ns; -- sim_handshake test
CONSTANT int_time   : TIME := 26500 ns + 0 * 40 ns;

-- Demoboard specific signals

SIGNAL leds_n       : UNSIGNED(3 DOWNTO 0);
SIGNAL keys_n       : UNSIGNED(3 DOWNTO 0);

BEGIN

-- ---------------------------------------------------------------------
-- demoboard pins
-- ---------------------------------------------------------------------

keys_n(0)          <= int_n;
keys_n(3 DOWNTO 1) <= (OTHERS => '0');

-- ---------------------------------------------------------------------
-- Test vector generation
-- ---------------------------------------------------------------------

int_n  <= '1', '0' AFTER int_time, '1' AFTER int_time + 600 ns;

bitout <= '1' WHEN  leds_n(0) = '0' OR (debug = '1' AND host_reg = 16#4002#)  ELSE '0';

-- ---------------------------------------------------------------------
-- Communicating with the uCore debugger via umbilical
-- ---------------------------------------------------------------------

make_initROM: IF  prog_len /= 0  GENERATE
   debug_mem: program_rom PORT MAP(debug_addr, debug_data);
END GENERATE make_initROM;

umbilical_proc: PROCESS

	VARIABLE text  : line;

   PROCEDURE tx_byte (number : IN byte) IS
   BEGIN
     WHILE  sending = '1' LOOP WAIT FOR cycle; END LOOP;
     send_byte <= '1';
     tx_buf <= number;
     WAIT UNTIL sending = '1';
     send_byte <= '0';
     tx_buf <= (OTHERS => 'Z');
   END tx_byte;

   PROCEDURE tx_word (number : IN data_bus) IS
   BEGIN
     out_buf <= (OTHERS => '0');
     out_buf(data_width-1 DOWNTO 0) <= number;
     FOR  i IN octetts DOWNTO 1  LOOP
        tx_byte(out_buf(i*8-1 DOWNTO (i-1)*8));
     END LOOP;
   END tx_word;

   PROCEDURE wait_ack IS
   BEGIN
      WHILE NOT (host_full = '1' AND host_buf = mark_ack) LOOP  WAIT FOR cycle;  END LOOP;
      WAIT UNTIL host_full = '0';
   END wait_ack;

   PROCEDURE rx_word (number : IN data_bus) IS
   BEGIN
      WHILE NOT (host_full = '1' AND host_reg(data_width-1 DOWNTO 0) = number)  LOOP  WAIT FOR cycle;  END LOOP;
      WAIT UNTIL host_full = '0';
   END rx_word;

   PROCEDURE rx_debug (number : IN data_bus) IS
   BEGIN
      WHILE NOT (host_full = '1' AND host_reg(data_width-1 DOWNTO 0) = number)  LOOP  WAIT FOR cycle;  END LOOP;
      host_ack <= '1';
      WAIT UNTIL host_full = '0';
      WAIT FOR cycle;
      host_ack <= '0';
   END rx_debug;

   PROCEDURE rx_byte (number : IN byte) IS
   BEGIN
      WHILE NOT (host_full = '1' AND host_reg(7 DOWNTO 0) = number)  LOOP  WAIT FOR cycle;  END LOOP;
      WAIT FOR cycle;
   END rx_byte;

   PROCEDURE tx_debug ( number : IN data_bus) IS
   BEGIN
      tx_byte(mark_debug);
      tx_word(number);
      wait_ack;
   END tx_debug;

BEGIN
--   switch_n     <= (OTHERS => '0');
   reset_n      <= '0';
   send_byte    <= '0';
   tx_buf       <= "ZZZZZZZZ";
   host_ack     <= '0';
   downloading  <= '0';
   uploading    <= '0';
   debug_addr   <= (OTHERS => '0');
   WAIT FOR 1000 ns;
   reset_n      <= '1';

   WAIT FOR 20 us;

   IF  prog_len /= 0 AND progload = '1'  THEN
		text := NEW string'("starting progload test ...");
      writeline(output, text);

-- send a string of NAK's, just in case
      FOR  i IN octetts DOWNTO 1  LOOP
         tx_byte(mark_nack);
      END LOOP;

-- load memory with reset
      tx_byte(mark_reset);  -- $CC
      tx_word(to_unsigned(0, data_width));        -- start address
      tx_word(to_unsigned(prog_len, data_width)); -- length
      FOR  i IN 0 TO  prog_len-1  LOOP         -- transfer memory image
         debug_addr <= to_unsigned(i, prog_addr_width);
         tx_byte(debug_data);
      END LOOP;
      wait_ack;
		text := NEW string'("progload test ok ");
      writeline(output, text);
      WAIT;
   END IF;

   IF  handshake = '1'  THEN -- debugger handshake see: monitor.fs
		text := NEW string'("starting handshake test ...");
      writeline(output, text);
      tx_debug(to_unsigned(0, data_width));
      rx_debug(slice('1', data_width));
      tx_debug(to_unsigned(16#3F5#, data_width));
      rx_debug(to_unsigned(16#305#, data_width));
      tx_debug(to_unsigned(0, data_width));
-- entering monitor loop
      rx_debug (to_unsigned(0, data_width)); -- now monitor waits for executable address

-- transfer "#c-bitout Ctrl-reg ! EXIT" to addr $200 and execute it
      tx_byte(mark_start);
      tx_word(to_unsigned(16#200#, data_width)); -- addr
      tx_word(to_unsigned( 6, data_width));      -- length
      tx_byte(to_unsigned(exp2(c_bitout) + 128, 8));
      tx_byte(op_NOOP);
      tx_byte(unsigned(to_signed(CTRL_REG, 8)));
      tx_byte(op_STORE);
      tx_byte(op_DROP);
      tx_byte(op_EXIT);
      wait_ack; -- now uCore waits for an execution address
      tx_debug(to_unsigned(16#200#, data_width)); -- execute it
      rx_debug (to_unsigned(0, data_width));
      tx_byte(mark_ack);
		text := NEW string'("handshake test ok ");
      writeline(output, text);
      WAIT;
   END IF;

   IF  debug = '1'  THEN
		text := NEW string'("starting debug register test ...");
      writeline(output, text);
      tx_debug(to_unsigned(16#8001#, data_width));
      rx_debug(to_unsigned(16#8001#, data_width));
      tx_debug(to_unsigned(16#4002#, data_width));
      rx_debug(to_unsigned(16#4002#, data_width));
      tx_byte(mark_ack);
      WHILE  sending = '1'  LOOP WAIT FOR baud/2;  END LOOP;
		text := NEW string'("debug register test ok ");
      writeline(output, text);
      WAIT;
   END IF;

   IF  upload = '1'  THEN  -- upload to data memory
		text := NEW string'("starting upload test ...");
      writeline(output, text);
      WAIT FOR 0 * 40 ns;
      uploading <= '1';
      tx_byte(mark_upload);
      IF  byte_addr_width = 0  THEN            -- cell addressing
         tx_word(to_unsigned( 8, data_width)); -- start address internal memory
         tx_word(to_unsigned( 4, data_width)); -- length
         FOR i IN 1 TO 4 LOOP
            tx_word(to_unsigned((16+i), data_width));
         END LOOP;
      ELSE                                     -- byte addressing
         tx_word(to_unsigned( 8 * bytes_per_cell, data_width)); -- start address internal memory
         tx_word(to_unsigned( 6, data_width)); -- length
         FOR i IN 1 TO 6 LOOP
            tx_byte(to_unsigned((16+i), 8));
         END LOOP;
      END IF;
      wait_ack;
      uploading <= '0';
      WAIT FOR cycle;
      IF  WITH_EXTMEM  THEN
         uploading <= '1';
         tx_byte(mark_upload);
         tx_word(to_unsigned(exp2(cache_addr_width), data_width)); -- start address external memory
         tx_word(to_unsigned( 4, data_width));                     -- length
         FOR i IN 5 TO 8 LOOP
            tx_word(to_unsigned((32+i), data_width));
         END LOOP;
         wait_ack;
         uploading <= '0';
      END IF;
      WHILE  bitout = '0'  LOOP WAIT FOR cycle;  END LOOP;
		text := NEW string'("upload test ok ");
      writeline(output, text);
      WAIT;
   END IF;

   IF  download = '1'  THEN  -- download from data memory
		text := NEW string'("starting download test ...");
      writeline(output, text);
      WAIT FOR 1200 ns + 3 * 40 ns;
      downloading <= '1';
      tx_byte(mark_download);
      tx_word(to_unsigned(bytes_per_cell, data_width));     -- start address internal memory
      tx_word(to_unsigned(8, data_width)); -- length
      IF  byte_addr_width = 0  THEN
         rx_word(to_unsigned(16#2211#, data_width));
         rx_word(to_unsigned(16#2211#, data_width));
         rx_word(to_unsigned(16#2211#, data_width));
         rx_word(to_unsigned(16#2211#, data_width));
         rx_word(to_unsigned(16#2211#, data_width));
         rx_word(to_unsigned(16#2211#, data_width));
         rx_word(to_unsigned(16#2211#, data_width));
         rx_word(to_unsigned(16#2211#, data_width));
         IF  WITH_EXTMEM  THEN
            tx_byte(mark_ack);
            WHILE  sending = '1'  LOOP WAIT FOR baud/2;  END LOOP;
            downloading <= '0';
            WAIT FOR baud;
            downloading <= '1';
            tx_byte(mark_download);
            tx_word(to_unsigned(exp2(cache_addr_width), data_width)); -- start address external memory
            tx_word(to_unsigned(2, data_width)); -- length
            rx_word(to_unsigned(16#6655#, data_width));
            rx_word(to_unsigned(16#8877#, data_width));
         END IF;
      ELSE
         rx_byte(to_unsigned(16#11#, 8));
         rx_byte(to_unsigned(16#22#, 8));
         rx_byte(to_unsigned(16#00#, 8));
         rx_byte(to_unsigned(16#00#, 8));
         rx_byte(to_unsigned(16#11#, 8));
         rx_byte(to_unsigned(16#22#, 8));
         rx_byte(to_unsigned(16#00#, 8));
         rx_byte(to_unsigned(16#00#, 8));
      END IF;
      tx_byte(mark_ack);
      WHILE  sending = '1'  LOOP WAIT FOR baud/2;  END LOOP;
      downloading <= '0';
		text := NEW string'("download test ok ");
      IF  bitout = '0'  THEN
         writeline(output, text);
      END IF;
      WAIT;
   END IF;

   IF  break = '1'  THEN -- multitasking: put terminal to sleep
		text := NEW string'("starting break test ...");
      writeline(output, text);
      WAIT FOR 80 us;
      tx_byte(mark_break);  -- put terminal to sleep
      WAIT FOR 80 us;
      tx_byte(mark_nbreak); -- wake terminal again
      WHILE  bitout = '0'  LOOP WAIT FOR cycle;  END LOOP;
		text := NEW string'("break test ok ");
      writeline(output, text);
      WAIT;
   END IF;

-- coretest
   text := NEW string'("starting core test ...");
   writeline(output, text);
   WAIT UNTIL bitout = '1';
   WAIT UNTIL bitout = '0';
   WAIT UNTIL bitout = '1';
   ASSERT false REPORT "core test ok" SEVERITY note;
   WAIT;

END PROCESS umbilical_proc;

to_target_proc: PROCESS
   VARIABLE number : byte := (OTHERS => 'Z');
BEGIN
   host_txd <= '1';
   sending <= '0';
   WAIT FOR 980 ns;
   LOOP
      WHILE  host_ack = '0' AND send_byte = '0'  LOOP  WAIT FOR cycle; END LOOP;
      sending <= '1';
      IF  host_ack = '1'  THEN
         number := mark_ack;
      ELSE
         number := tx_buf;
      END IF;
      host_txd <= '0';  -- start bit
      WAIT FOR baud;
      FOR  i IN 0 TO 7  LOOP
        host_txd <= number(i);
        WAIT FOR baud;
      END LOOP;
      host_txd <= '1';  -- stop bit
      sending <= '0';
      WAIT FOR baud;   -- wait for full stop bit
   END LOOP;
END PROCESS to_target_proc ;

from_target_proc : PROCESS

   PROCEDURE rx_uart IS
   BEGIN
     WHILE  host_rxd /= '0'  LOOP WAIT FOR cycle/2; END LOOP;
     WAIT FOR baud/2;
     FOR  i IN 0 TO 7  LOOP
        WAIT FOR baud;
        host_buf(i) <= host_rxd;
     END LOOP;
     WAIT FOR baud/2;
   END rx_uart;

BEGIN
   host_full <= '0';
   host_reg <= (OTHERS => '1');
   WAIT FOR 1 us;
   LOOP
      WAIT FOR cycle;
      host_full <= '0';
      WHILE  host_rxd = '1'  LOOP WAIT FOR cycle;  END LOOP;
      IF  downloading = '1'  THEN
         IF  byte_addr_width = 0  THEN
            FOR i IN octetts-1 DOWNTO 0 LOOP
               rx_uart;
               host_reg <= host_reg(host_reg'high-8 DOWNTO 0) & host_buf;
            END LOOP;
         ELSE
            rx_uart;
            host_reg <= resize(host_buf, host_reg'length);
         END IF;
         host_full <= '1';
      ELSE
         rx_uart;
         IF  host_buf = mark_ack  THEN
            host_full <= '1';
         ELSIF  host_buf = mark_debug  THEN
            FOR i IN octetts-1 DOWNTO 0 LOOP
               rx_uart;
               host_reg <= host_reg(host_reg'high-8 DOWNTO 0) & host_buf;
            END LOOP;
            host_full <= '1';
         END IF;
      END IF;
   END LOOP;

END PROCESS from_target_proc ;

-- ---------------------------------------------------------------------
-- The clock oscillator
-- ---------------------------------------------------------------------

xtal_clock: PROCESS
BEGIN
  xtal <= '0';
  WAIT FOR 500 ns;
  LOOP
    xtal <= '1';
    WAIT FOR xtal_cycle/2;
    xtal <= '0';
    WAIT FOR xtal_cycle/2;
  END LOOP;
END PROCESS xtal_clock;

-- ---------------------------------------------------------------------
-- external SDRAM
-- ---------------------------------------------------------------------

-- ---------------------------------------------------------------------
-- uCore FPGA
-- ---------------------------------------------------------------------

myFPGA: fpga PORT MAP (
   reset_n    => reset_n,
   clock      => xtal,
-- Demoboard specific pins                    
   keys_n     => keys_n,
--   beep       => OUT   STD_LOGIC;
   leds_n     => leds_n,
-- temp sensor
--   SCL        => OUT   STD_LOGIC;
--   SDA        => INOUT STD_LOGIC;
-- serial E2prom
--   I2C_SCL    => OUT   STD_LOGIC;
--   I2C_SDA    => INOUT STD_LOGIC;
-- IR es ist mir unklar, ob das ein Sender oder ein Empf�nger ist, deshal erstmal auskommentiert
--   IR         => ????? STD_LOGIC;
-- VGA
--   VGA_HSYNC  => OUT   STD_LOGIC;
--   VGA_VSYNC  => OUT   STD_LOGIC;
--   VGA_BGR    => OUT   UNSIGNED(2 DOWNTO 0);
-- LCD                                        
--   LCD_RS     => OUT   STD_LOGIC;
--   LCD_RW     => OUT   STD_LOGIC;
--   LCD_E      => OUT   STD_LOGIC;
--   LCD_Data   => OUT   UNSIGNED(7 DOWNTO 0);
-- 7-Segment                                  
--   DIG        => OUT   UNSIGNED(3 DOWNTO 0);
--   SEG        => OUT   UNSIGNED(7 DOWNTO 0);
-- SDRAM                                      
--   SD_DQ      => INOUT UNSIGNED(15 DOWNTO 0);
--   SD_A       => OUT   UNSIGNED(11 DOWNTO 0);
--   SD_BA      => OUT   UNSIGNED( 1 DOWNTO 0);
--   SD_LDQM    => OUT   STD_LOGIC;
--   SD_UDQM    => OUT   STD_LOGIC;
--   SD_CKE     => OUT   STD_LOGIC;
--   SD_CLK     => OUT   STD_LOGIC;
--   SD_CS_n    => OUT   STD_LOGIC;
--   SD_RAS_n   => OUT   STD_LOGIC;
--   SD_CAS_n   => OUT   STD_LOGIC;
--   SD_WE_n    => OUT   STD_LOGIC;
-- umbilical port for debugging
   dsu_rxd    => host_txd, -- host -> target
   dsu_txd    => host_rxd  -- target -> host
);

END testbench;
